package observer_real_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "observer_real_util.svh"
endpackage : observer_real_pkg