package manipulator_strg_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "manipulator_strg_util.svh"
endpackage : manipulator_strg_pkg